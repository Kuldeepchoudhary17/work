magic
tech sky130A
timestamp 1637227170
<< nmos >>
rect 200 -260 300 0
<< ndiff >>
rect 0 -20 200 0
rect 0 -240 20 -20
rect 180 -240 200 -20
rect 0 -260 200 -240
rect 300 -20 500 0
rect 300 -240 320 -20
rect 480 -240 500 -20
rect 300 -260 500 -240
<< ndiffc >>
rect 20 -240 180 -20
rect 320 -240 480 -20
<< poly >>
rect 200 0 300 18
rect 200 -278 300 -260
<< locali >>
rect 10 -20 190 -10
rect 10 -240 20 -20
rect 180 -240 190 -20
rect 10 -250 190 -240
rect 310 -20 490 -10
rect 310 -240 320 -20
rect 480 -240 490 -20
rect 310 -250 490 -240
<< end >>
