* SPICE3 file created from nmos.ext - technology: sky130A

X0 a_300_n260# a_200_n278# a_0_n260# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.6e+06u l=1e+06u
