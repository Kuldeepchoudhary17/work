magic
tech sky130A
timestamp 1637226432
<< nwell >>
rect -18 -518 518 18
<< pmos >>
rect 200 -500 300 0
<< pdiff >>
rect 0 -20 200 0
rect 0 -480 20 -20
rect 180 -480 200 -20
rect 0 -500 200 -480
rect 300 -20 500 0
rect 300 -480 320 -20
rect 480 -480 500 -20
rect 300 -500 500 -480
<< pdiffc >>
rect 20 -480 180 -20
rect 320 -480 480 -20
<< poly >>
rect 200 0 300 18
rect 200 -518 300 -500
<< locali >>
rect 10 -20 190 -10
rect 10 -480 20 -20
rect 180 -480 190 -20
rect 10 -490 190 -480
rect 310 -20 490 -10
rect 310 -480 320 -20
rect 480 -480 490 -20
rect 310 -490 490 -480
<< end >>
